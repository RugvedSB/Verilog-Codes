`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Name : Rugved Bopardikar
// 
// Design Name: Full Adder
// Module Name: full_adder
// Project Name: 
// Target Devices: Basys 3 Artix 7
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module half_adder(
    input wire a, b,
    output sout,
    output cout
    );
    
assign sout = a ^ b;
assign cout = a & b;

endmodule

module full_adder(
    input a, b, cin,
    output s,
    output c
    );
    
wire t1, t2, t3;

half_adder h1(a, b, t1, t2);
half_adder h2(t1, cin, s, t3);

assign c = t2 | t3;

endmodule 